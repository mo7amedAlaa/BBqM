module FSM ( clk , reset , pCount , switch1 , switch2 , con ) ;
       input clk , reset , switch1 , switch2 ;
       input  [2:0] pCount;
       output [4:0] con;

       parameter S0 = 2'b00 ,
                 S1 = 2'b01 , 
                 S2 = 2'b10 ,
					  S3 = 2'b11 ;

       reg [1:0] tCount ;

       always @(*)
       begin
           if(reset) 
             begin
               tCount = S0 ;
             end
           else
             begin
                   if( ~switch1 && switch2 )
                           tCount <= S1 ;
                    else if( switch1 && ~switch2 )
                           tCount <= S2 ;                   
                    else if( switch1 && switch2 )
                           tCount <= S3 ;
             end
        end

      assign con = { tCount , pCount } ;

endmodule

module decoder_7seg (A, B, C, D, led_a, led_b, led_c, led_d, led_e, led_f, led_g);
 
 input A, B, C, D; 
 output led_a, led_b, led_c, led_d, led_e, led_f, led_g;

  assign led_a = ~(A | C | B&D | ~B&~D); 
  assign led_b = ~(~B | ~C&~D | C&D);
  assign led_c = ~(B | ~C | D); 
  assign led_d = ~(~B&~D | C&~D | B&~C&D | ~B&C |A); 
  assign led_e = ~(~B&~D | C&~D);
  assign led_f = ~(A | ~C&~D | B&~C | B&~D); 
  assign led_g = ~(A | B&~C | ~B&C | C&~D); 
 
endmodule

